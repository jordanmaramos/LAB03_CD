library verilog;
use verilog.vl_types.all;
entity MUX_4X1_vlg_vec_tst is
end MUX_4X1_vlg_vec_tst;
