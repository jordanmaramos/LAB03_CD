library verilog;
use verilog.vl_types.all;
entity LAB03_vlg_check_tst is
    port(
        MUX_OUT         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end LAB03_vlg_check_tst;
