library verilog;
use verilog.vl_types.all;
entity MUX_2X1_COMPORT_vlg_vec_tst is
end MUX_2X1_COMPORT_vlg_vec_tst;
