library verilog;
use verilog.vl_types.all;
entity MUX_2X1_LOGIC_vlg_check_tst is
    port(
        D               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MUX_2X1_LOGIC_vlg_check_tst;
