library verilog;
use verilog.vl_types.all;
entity MUX_4X1_vlg_check_tst is
    port(
        D               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MUX_4X1_vlg_check_tst;
