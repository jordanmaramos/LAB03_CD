library verilog;
use verilog.vl_types.all;
entity MUX_2X1_LOGIC_vlg_vec_tst is
end MUX_2X1_LOGIC_vlg_vec_tst;
