library verilog;
use verilog.vl_types.all;
entity LAB03 is
    port(
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        A3              : in     vl_logic;
        B0              : in     vl_logic;
        B1              : in     vl_logic;
        MUX_OUT         : out    vl_logic
    );
end LAB03;
